 	//THIS IS GENERATED FILE!
	parameter ROM0_DATA='h4b1;
	parameter ROM_PATH="/home/ic_contest/509/CRYSTALS/HDL";
