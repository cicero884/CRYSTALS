/********
define MUL_STAGE_CNT for controller to control out_en and clk gating
change depend on your design of mo_mul
********/
`define MUL_STAGE_CNT `DATA_WIDTH
