module butterfly (
	
)
