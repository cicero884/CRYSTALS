 	`define ROM0_DATA 'h4b1
	`define ROM_PATH "/home/cicero/code/CRYSTALS/HDL" 
