module ntt (
	input clk,input reset,
	input in_en,input data_in,
	output logic addr,output logic data_out,
	output logic done
);
always

endmodule
