// if you change to your mo_mul
// you dont need to include ntt.svh
// just change MUL_STAGE_CNT to your design
`include "ntt.svh"
`define MUL_STAGE_CNT `DATA_WIDTH
