/**********
change depend on add_sub design
**********/
`ifndef ADD_SUB_SVH
`define ADD_SUB_SVH

`define ADD_SUB_STAGE_CNT 2

`endif
