// convert macro value to string
`define STRINGIFY(x) `"x`"
