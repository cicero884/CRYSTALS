 	//THIS IS GENERATED FILE!
	`define MULTYPE_KRED
