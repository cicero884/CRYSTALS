/**********
change depend on add_sub design
**********/
parameter ADD_SUB_STAGE_CNT=2;
