/**********
change depend on add_sub design
**********/
parameter NTT_ADD_SUB_STAGE_CNT =1;
parameter INTT_ADD_SUB_STAGE_CNT=2;
