`define ADD_SUB_STAGE_CNT 2
