 	`define Q 3329
	`define NTT_STAGE_CNT 7 
